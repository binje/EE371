module divider8 (quotient, remainder, op1, op2);
	parameter WIDTH = 8;
	output [(WIDTH-1):0] out, remainder;
	input [(WIDTH-1):0] op1, op2;
	
	
endmodule 