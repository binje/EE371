module alu (out, func, op1, op2);
	input [1:0] func;
	input [7:0] op1, op2;
	output [7:0] out;
	
endmodule 