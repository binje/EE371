library verilog;
use verilog.vl_types.all;
entity recognize6_testbench is
end recognize6_testbench;
