module syncDown (clk)