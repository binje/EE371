library verilog;
use verilog.vl_types.all;
entity recognize3_testbench is
end recognize3_testbench;
